module dand(input a, input b, output c);
	assign #1 c = a && b;
endmodule