module XOR1(input xin0, input xin1, output wire xout);
	assign xout = xin0 ^ xin1;
endmodule