module top(input in0, input in1, input in2, input[1:0] in3, output wire[6:0] out);
	wire cout;
	wire sum;
	wire par;
	wire muxout;
	wire[1:0] compout;
	
	sumator DUT1(.cin(in0),.in0(in1),.in1(in2),.cout(cout),.par(par),.sum(sum));
	comparatort DUT2(.in0(in3),.in1(1'h1),.out(compout));
	muxt DUT3(.in2(cout),.in0(sum),.in1(par),.sel(compout),.out(muxout));
	transcodor DUT4(.in(muxout),.out(out));
endmodule