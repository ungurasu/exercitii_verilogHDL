module parityChecker(input in, output wire out);
	assign out = !in;
endmodule