module bancadetestare();
	reg[2:0] a;
	reg[2:0] b;
	reg[2:0] c;
	reg[2:0] d;
	reg[2:0] e;
	reg[2:0] opcode;
	reg sel_1;
	reg[1:0] sel_2;
	wire[2:0] out;
	wire carry_out;
	
	toptema DUT1(.a(a), .b(b), .c(c), .d(d), .e(e), .opcode(opcode), .sel_1(sel_1), .sel_2(sel_2), .out(out), .carry_out(carry_out));	
	initial begin
		sel_1 = 0;
		sel_2 = 0;
		opcode = 0;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 0;
		opcode = 1;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 0;
		opcode = 2;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 0;
		opcode = 3;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 0;
		opcode = 4;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 0;
		opcode = 5;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 1;
		opcode = 0;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 2;
		opcode = 0;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 1;
		sel_2 = 2;
		opcode = 0;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
		sel_1 = 0;
		sel_2 = 3;
		opcode = 0;
		a = 2;
		b = 3;
		c = 2;
		d = 3;
		e = 2;
		#20;
	end
endmodule