`timescale 1ns/1ps

module testbench();
	reg[3:0] addr;
	reg[3:0] addrop1;
	reg[3:0] addrop2;
	reg[3:0] data;
	reg clock;
	reg we;
	reg sel;
	reg[1:0] opcode;
	wire[4:0] out;
	
	TOPt DUT1(.clock(clock),.addr(addr),.addrop1(addrop1),.addrop2(addrop2),.data(data),.we(we),.opcode(opcode),.sel(sel),.out(out));
	
	initial begin
		clock <= 1;
		repeat (33) 
			#21 clock <= !clock;
	end
	
	initial begin
		we = 0;
		sel = 0;
		#42;
		addr = 0;
		data = 10;
		we = 1;
		sel = 0;
		#42;
		addr = 1;
		data = 12;
		we = 1;
		sel = 0;
		#42;
		addr = 2;
		data = 5;
		we = 1;
		sel = 0;
		#42;
		addr = 3;
		data = 6;
		we = 1;
		sel = 0;
		#42;
		addr = 4;
		data = 14;
		we = 1;
		sel = 0;
		#42;
		addr = 5;
		data = 20;
		we = 1;
		sel = 0;
		#42;
		addr = 6;
		data = 15;
		we = 0;
		sel = 0;
		#42;
		addr = 6;
		data = 15;
		we = 0;
		sel = 0;
		addrop1 = 0;
		addrop2 = 4;
		opcode = 0;
		#42;
		addr = 6;
		data = 15;
		we = 0;
		sel = 0;
		addrop1 = 2;
		addrop2 = 2;
		opcode = 1;
		#42;
		addr = 6;
		data = 15;
		we = 0;
		sel = 0;
		addrop1 = 4;
		addrop2 = 1;
		opcode = 2;
		#42;
		addr = 6;
		data = 15;
		we = 0;
		sel = 0;
		addrop1 = 1;
		addrop2 = 5;
		opcode = 3;
		#42;
		addr = 6;
		data = 15;
		we = 0;
		sel = 1;
		addrop1 = 0;
		addrop2 = 2;
		opcode = 3;
		#42;
		addr = 3;
		data = 15;
		we = 0;
		sel = 1;
		addrop1 = 6;
		addrop2 = 3;
		opcode = 3;
		#42;
		addr = 2;
		data = 15;
		we = 0;
		sel = 1;
		addrop1 = 6;
		addrop2 = 3;
		opcode = 3;
		#42;
		addr = 3;
		data = 15;
		we = 0;
		sel = 1;
		addrop1 = 6;
		addrop2 = 3;
		opcode = 3;
		#42;
		addr = 4;
		data = 15;
		we = 0;
		sel = 1;
		addrop1 = 6;
		addrop2 = 3;
		opcode = 3;
		#42;
		addr = 5;
		data = 15;
		we = 0;
		sel = 1;
		addrop1 = 6;
		addrop2 = 3;
		opcode = 3;
		#42;
	end
endmodule